`include "alu.v"
`include "alu_control.v"
`include "control.v"
`include "im.v"
`include "mux2.v"
`include "registers.v"

module single_cycle ();

    

endmodule // single_cycle
